----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:19:45 04/21/2011 
-- Design Name: 
-- Module Name:    FILE_SELECT_FIXE - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FILE_SELECT_FIXE is
    Port ( FILE_SELECT : out  STD_LOGIC_VECTOR (7 downto 0));
end FILE_SELECT_FIXE;

architecture Behavioral of FILE_SELECT_FIXE is

begin
FILE_SELECT<="00010000";

end Behavioral;

