-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity AZRAEL_256x256_ROM is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of AZRAEL_256x256_ROM is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_01 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_02 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_03 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_04 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_05 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_09 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_11 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_12 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_13 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_14 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_15 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_16 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_17 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_18 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_19 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_20 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_21 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_22 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_24 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_25 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_26 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_27 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_28 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_31 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_35 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_36 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_37 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_38 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFF003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_04 of inst : label is "FFFFFFFFFE7FF8000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFE3FC00000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFF";
    attribute INIT_06 of inst : label is "FFFFFFFFFF00000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFF";
    attribute INIT_07 of inst : label is "FFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFF";
    attribute INIT_08 of inst : label is "FFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000007FFFFF";
    attribute INIT_09 of inst : label is "FFFFFFFFFE2000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_0A of inst : label is "FFFFFFFFFE2000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_0B of inst : label is "FFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_0C of inst : label is "FFFFFFFFFF00000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFF0000007FFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFF04000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFF80000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFE0000007FFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFC0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF80000007FFFFF";
    attribute INIT_11 of inst : label is "FFFFFFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFF00000007FFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFE60000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFC00000007FFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFE70000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF80000000FFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFE30000000000000FFFFFFFFFFFFFFFFFFFFFFFFFE000000007FFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFF38000000000000FFFFFFFFFFFFFFFFFFFFFFFFF800000000FFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFF18000000000000FFFFFFFFFFFFFFFFFFFFFFFFE000000001FFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFF8C000000000000FFFFFFFFFFFFFFFFFFFFFFFFC000000003FFFFFF";
    attribute INIT_18 of inst : label is "FFFFFFFFFF88000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000007FFFFFF";
    attribute INIT_19 of inst : label is "FFFFFFFFFFC0000000000000FFFFFFFFFFFFFFFFFFFFFFFC000000000FFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFF9C0000000000000FFFFFFFFFFFFFFFFFFFFFFF0000000000FFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFF9C0000000000000FFFFFFFFFFFFFFFFFFFFFFC0000000001FFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFF9C0000000000000FFFFFFFFFFFFFFFFFFFFFF00000000001FFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFCC0000000000000FFFFFFFFFFFFFFFFFFFFFC00000000003FFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFEC00000000000007FFFFFFFFFFFFFFFFFFFF000000000007FFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFE400007FF8000003FFFFFFFFFFFFFFFFFFFC00000000000FFFFFFFF";
    attribute INIT_20 of inst : label is "FFFFFFFFFE00007FFF8000001FFFFFFFFFFFFFFFFFFF000000000001FFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFE000003FF80000003FFFFFFFFFFFFFFFFF8000000000007FFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFE0000007F00000001FFFFFFFFFFFFFFFFF000000000000FFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFF800000007800000003FFFFFFFFFFFFFFF8000000000001FFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFF000000000000000000FFFFFFFFFFFFFFE0000000000003FFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFE0000000000000000003FFFFFFFFFFFFF80000000000007FFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFC00000000000000000003FFFFFFFFFFFE0000000000001FFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF800000000000000000000FFFFFFFFFFF00000000000003FFFFFFFFFF";
    attribute INIT_28 of inst : label is "FFFFFFFF80000000000000000000007FFFFFFFFC0000000000000FFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFF000000000000000000000003FFFFFFE00000000000001FFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFE0000000000000000000000003FFFFFC00000000000007FFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFE00000000000000000000000001FFFE00000000000001FFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFE000000000000000000000000003FF800000000000003FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFF8000000000000000000000000001E00000000000000FFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFC0000000000000000000000000000000000000000003FFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF80000000000000000000000000000000000000000007FFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "FFFFFFFC000000000000000000000000000000000000000001FFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "FFFFFFFE000000000000000000000000000000000000000007FFFFFFFFFFFFFF";
    attribute INIT_32 of inst : label is "FFFFFFFF00000000000000000000000000000000000000000FFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFF80000000000000000000000000000000000000003FFFFFFFFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFFC0000000000000000000000000000000000000007FFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFC000000000003000000000000000000000000001FFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFA000000000001800000000000000000000000007FFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFF3000000000001C0000000000000000000000000FFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFF180000000000020000000000000000000000003FFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFD18000000000000000000000000000000000000FFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFF988000000000000000000000000000000000003FFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFF8C4000000000000000000000000000000000007FFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFCC200004000000000000000000000000000001FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFC620001FF80000000000000000000000000007FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFE600003FFC000000000000000000000000000FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFE300003FFC000000000000000000000000003FFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0800067FFFFF";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8800067FFFFF";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8000047FFFFF";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFF007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C00007FFFFF";
    attribute INIT_04 of inst : label is "FFFFFFFFFE7FFC000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C00007FFFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFE3F80000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C00047FFFFF";
    attribute INIT_06 of inst : label is "FFFFFFFFFF08000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C00047FFFFF";
    attribute INIT_07 of inst : label is "FFFFFFFFFF800000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF88800C7FFFFF";
    attribute INIT_08 of inst : label is "FFFFFFFFFF80007FFC0001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8800067FFFFF";
    attribute INIT_09 of inst : label is "FFFFFFFFFE203F7FFC00007FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8C00067FFFFF";
    attribute INIT_0A of inst : label is "FFFFFFFFFE203C7978CFC03FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8E00047FFFFF";
    attribute INIT_0B of inst : label is "FFFFFFFFFE001F3000FFF80FFFFFFFFFFFFFFFFFFFFFFFFFFFFF8908047FFFFF";
    attribute INIT_0C of inst : label is "FFFFFFFFFE000F80000F7C07FFFFFFFFFFFFFFFFFFFFFFFFFFFF0018047FFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFF0C018000000F03FFFFFFFFFFFFFFFFFFFFFFFFFFFF0010047FFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFF8400800003C7C3FFFFFFFFFFFFFFFFFFFFFFFFFFFE14000C7FFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFC03600001703E1FFFFFFFFFFFFFFFFFFFFFFFFFFFE36008C7FFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFC0300000100731FFFFFFFFFFFFFFFFFFFFFFFFFFFC3800087FFFFF";
    attribute INIT_11 of inst : label is "FFFFFFFFFFE0380000000018FFFFFFFFFFFFFFFFFFFFFFFFFFF03800007FFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFE60198000000018FFFFFFFFFFFFFFFFFFFFFFFFFFE08800507FFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFE700180000020F0FFFFFFFFFFFFFFFFFFFFFFFFFFC38800C1FFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFE300EE000600360FFFFFFFFFFFFFFFFFFFFFFFFFE038000C0FFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFF3800C010000378FFFFFFFFFFFFFFFFFFFFFFFFFC0E000040FFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFF1C030710070030FFFFFFFFFFFFFFFFFFFFFFFFF01C000603FFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFF8C03C012070020FFFFFFFFFFFFFFFFFFFFFFFFC079010787FFFFFF";
    attribute INIT_18 of inst : label is "FFFFFFFFFF8C00F8138200B0FFFFFFFFFFFFFFFFFFFFFFFF00E261B38FFFFFFF";
    attribute INIT_19 of inst : label is "FFFFFFFFFFC01007F1E000C0FFFFFFFFFFFFFFFFFFFFFFFC000001238FFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFF9C00187F06038C0FFFFFFFFFFFFFFFFFFFFFFF81C0000071FFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFF9C003CC7C437850FFFFFFFFFFFFFFFFFFFFFFC0619C00061FFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFF9C02C000000E010FFFFFFFFFFFFFFFFFFFFFF00E38C083C3FFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFCC07C0000018010FFFFFFFFFFFFFFFFFFFFFC0020C00C787FFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFEC1C00000000000FFFFFFFFFFFFFFFFFFFFF00100E01B40FFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFE44000FFF8002203FFFFFFFFFFFFFFFFFFFC0180C6401C1FFFFFFFF";
    attribute INIT_20 of inst : label is "FFFFFFFFFE00007FFF85005C1FFFFFFFFFFFFFFFFFFF0000230E81C3FFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFE000007FF87C05407FFFFFFFFFFFFFFFFFC010030030007FFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFE000000FF84851601FFFFFFFFFFFFFFFFF007C07083E20FFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFF8000000078A8957003FFFFFFFFFFFFFFF800FE0039F6C1FFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFF0000000001A8051800FFFFFFFFFFFFFFE0019F0033EE07FFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFE007F3FC001FF0E16003FFFFFFFFFFFFF800F1F0003380FFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFC06D01FF000170803C003FFFFFFFFFFFE003F28000C381FFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF81F800C7F000300806000FFFFFFFFFFF00078381E00007FFFFFFFFFF";
    attribute INIT_28 of inst : label is "FFFFFFFF8E00000FF9801C0400F0007FFFFFFFFC0001470E471C0FFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFBC10000009C00400707C0003FFFFFFE0000000000F383FFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFE3E10000000600600380F00003FFFFFC000F8001838E07FFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFE0C100000C01C0600C1C3F00001FFFE000EFC00183B81FFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFE07000000807C030100003800007FF8000E000181B003FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFF87800000003003013FC018C00003C001EF002000780FFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFF801800000403607600000000000000001C0806038E03FFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF820800004001C06E0000008178000000000000031C07FFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "FFFFFFFC0080801F001E068800001C3FE0000000000E006703FFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "FFFFFFFE00088000C10006600000002007000000000E070407FFFFFFFFFFFFFF";
    attribute INIT_32 of inst : label is "FFFFFFFF00300000C100092000000200000003000006FF880FFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFF80300F01800001C0003826E000C01800000071C03FFFFFFFFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFFC00600F30018018000FC06E00000100000007F00FFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFC00200FC0070308002C7020000C7000000000C03FFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFE060FF7800701C000E830020018607000001F807FFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFF30F1007120421C000E3018388C0000800003E01FFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFF389800005006070022781800E00000606007007FFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFD1C0000001C00000000000000C0000000001E00FFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFF98C6000000CB18000000000000000FE0181F803FFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFF8C670000003B1C0000000000800000018E7180FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFCC660004003004000000000000000000820981FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFC620223FF82207800000000400000038000E07FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFE600783FFC0203C000001F040000007809880FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFE301703FFC02005EFF9FCFE00000002028E03FFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF";
    attribute INIT_01 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFF";
    attribute INIT_02 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_03 of inst : label is "FFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_04 of inst : label is "FFFFFFFFFE7FFC000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_05 of inst : label is "FFFFFFFFFE3FE0000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_06 of inst : label is "FFFFFFFFFF1C000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_07 of inst : label is "FFFFFFFFFF8003FFFF0007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_08 of inst : label is "FFFFFFFFFF801FFFFFFC01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFF";
    attribute INIT_09 of inst : label is "FFFFFFFFFE60FFFFFFFFE07FFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF7FFFFF";
    attribute INIT_0A of inst : label is "FFFFFFFFFE20FFFFFFFFF83FFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF7FFFFF";
    attribute INIT_0B of inst : label is "FFFFFFFFFE307FFFFFFFFE0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF7FFFFF";
    attribute INIT_0C of inst : label is "FFFFFFFFFE1C3FFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFF7FFFFF";
    attribute INIT_0D of inst : label is "FFFFFFFFFF0E7FFFFFFFFFC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFF7FFFFF";
    attribute INIT_0E of inst : label is "FFFFFFFFFF8FFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFFF7FFFFF";
    attribute INIT_0F of inst : label is "FFFFFFFFFFC7FFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFF7FFFFF";
    attribute INIT_10 of inst : label is "FFFFFFFFFFC3FFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFE7FFFFF";
    attribute INIT_11 of inst : label is "FFFFFFFFFFE1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9FFFFFC7FFFFF";
    attribute INIT_12 of inst : label is "FFFFFFFFFE707FFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFF";
    attribute INIT_13 of inst : label is "FFFFFFFFFE703FFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFC7FFFFF9FFFFFF";
    attribute INIT_14 of inst : label is "FFFFFFFFFE383FFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFF0FFFFFF";
    attribute INIT_15 of inst : label is "FFFFFFFFFF3E1FFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFF1FFFFFF";
    attribute INIT_16 of inst : label is "FFFFFFFFFF3F9FFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFF1FFFFFFC7FFFFFF";
    attribute INIT_17 of inst : label is "FFFFFFFFFF9DFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFEFFFFFFF";
    attribute INIT_18 of inst : label is "FFFFFFFFFF8DFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFEFFFFFFF";
    attribute INIT_19 of inst : label is "FFFFFFFFFFCDFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFE1FFFFFFFFFFFFFFF";
    attribute INIT_1A of inst : label is "FFFFFFFFFDC1FFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFBFFFFFFF";
    attribute INIT_1B of inst : label is "FFFFFFFFF9C1FFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFE0FFFFFFFF1FFFFFFF";
    attribute INIT_1C of inst : label is "FFFFFFFFFDC1FFE00043FFF9FFFFFFFFFFFFFFFFFFFFFF83FFFFFFFF3FFFFFFF";
    attribute INIT_1D of inst : label is "FFFFFFFFFCE1FF000003FFF8FFFFFFFFFFFFFFFFFFFFFE0FFFFFFFFC7FFFFFFF";
    attribute INIT_1E of inst : label is "FFFFFFFFFEEFFF00FF83FFFCFFFFFFFFFFFFFFFFFFFFF83FFFFFFFFDFFFFFFFF";
    attribute INIT_1F of inst : label is "FFFFFFFFFE47FEFFFF87FFFC7FFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFF";
    attribute INIT_20 of inst : label is "FFFFFFFFFE0DF8FFFF8FFFFE1FFFFFFFFFFFFFFFFFFF03FFFFFFFFE7FFFFFFFF";
    attribute INIT_21 of inst : label is "FFFFFFFFFF00007FFF9FFFFF0FFFFFFFFFFFFFFFFFFC07FFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFE000001FF9FFFFF03FFFFFFFFFFFFFFFFF01FFFFFFFFFDFFFFFFFFF";
    attribute INIT_23 of inst : label is "FFFFFFFFF800FC000FDFFFFFC07FFFFFFFFFFFFFFFC03FFFFFFFFF3FFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFF80FFFF0031FFFFFF01FFFFFFFFFFFFFFF00FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFE0FFFFFF801FFFFFFE07FFFFFFFFFFFFF807FFFFFFFFF9FFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFE3FFFFFFF807FFFFFF807FFFFFFFFFFFE01FFFFFFFFFE3FFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFFC7FFFFFFFF83FFFFFFE01FFFFFFFFFFF807FFFFFFFFFCFFFFFFFFFFF";
    attribute INIT_28 of inst : label is "FFFFFFFFFFFFFFFFFFE0FFFFFFFC007FFFFFFFFC01FFFFFFFFFE1FFFFFFFFFFF";
    attribute INIT_29 of inst : label is "FFFFFFFFFFFFFFFFFFF87FFFFFFF0003FFFFFFF007FFFFFFFFFE7FFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFFFFFE7FFFFFFFFFFE3FFFFFFFE0003FFFFFC01FFFFFFFFFF8FFFFFFFFFFFF";
    attribute INIT_2B of inst : label is "FFFFFFFE3FFFFFFFFFFF1FFFFFFFFE0003FFFE007FFFFFFFFFC3FFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FFFFFFFF1FFFFFFFFFFF9FFFFFFFFFC0007FF801FFFFFFFFFF87FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFF8FFFFFFFFFFFDFFFFFFFFFF00003E007FFFFFFFFFE1FFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFF837FFFFFFFFFF8FFFFFC0FFFE0000001FFFFFFFFFFC7FFFFFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFF827FFFFFFFFFF8FFF8000FFFFF000007FFFFFFFFFF8FFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "FFFFFFFC03FFFFFFFFFF9FFE0007FFFFFFC003FFFFFFFFFFC3FFFFFFFFFFFFFF";
    attribute INIT_31 of inst : label is "FFFFFFFE03FFFFFFFFFF1FFC001FFFFFFFE00FFFFFFFFFFF8FFFFFFFFFFFFFFF";
    attribute INIT_32 of inst : label is "FFFFFFFF01FFFFFFFFFF1FF0007FFFFC0FE03FFFFFFFFFFC1FFFFFFFFFFFFFFF";
    attribute INIT_33 of inst : label is "FFFFFFFF80FFFFFFFFFF7FE001FFFFF80FFFFFFFFFFFFFF87FFFFFFFFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFFC0FFFFFFFFFF7FE007FFFFF80FFFFFFFFFFFFFF0FFFFFFFFFFFFFFFF";
    attribute INIT_35 of inst : label is "FFFFFFFFE2FFFFFFFFFF78C01FFFFFF81FFFFFFFFFFFFF83FFFFFFFFFFFFFFFF";
    attribute INIT_36 of inst : label is "FFFFFFFFF3FFFFFFFFFF7E003FFFFFFFFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFF";
    attribute INIT_37 of inst : label is "FFFFFFFF3FFFFFFFFFFF3E007FFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFF";
    attribute INIT_38 of inst : label is "FFFFFFFF3DFFFFFFFFFF9F00FFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFF";
    attribute INIT_39 of inst : label is "FFFFFFFD1DFFF00FFFFFC301FFFFFFFFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFF";
    attribute INIT_3A of inst : label is "FFFFFFF98DFE0000FFFFC003FFFFFFFFFFFFFFFFFFFF83FFFFFFFFFFFFFFFFFF";
    attribute INIT_3B of inst : label is "FFFFFFF8CEFE20001FFFF00001FF7FFFFFFFFFFFFFFE0FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFF8C6FFF3E00FFFFE000001FFFFFFFFFFFFFFFC3FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFC667FFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFF07FFFFFFFFFFFFFFFFFFF";
    attribute INIT_3E of inst : label is "FFFFFFFE713FFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3F of inst : label is "FFFFFFFE31BFF3FFE7FFFFFFFFFFFFFFFFFFFFFFFF87FFFFFFFFFFFFFFFFFFFF";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
