----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:59:34 12/21/2010 
-- Design Name: 
-- Module Name:    testdowntojeterpoubelle - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity testdowntojeterpoubelle is
    Port ( aa : in  STD_LOGIC_VECTOR (0 downto 7);
           zz : in  STD_LOGIC_VECTOR (7 downto 0));
end testdowntojeterpoubelle;

architecture Behavioral of testdowntojeterpoubelle is

begin


end Behavioral;

